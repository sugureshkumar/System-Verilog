class axi_gen;
	task run();
		$display("axi_gen:: run");
	endtask
endclass
