class abc;
	rand  int unsigned  a;

	constraint c1 {a inside{[0:9]};}	
	
endclass
