`include "axi_bfm.sv"
`include "axi_gen.sv"
`include "axi_cov.sv"
`include "axi_mon.sv"
`include "axi_env.sv"
`include "axi_tb.sv"
`include "top.sv"
