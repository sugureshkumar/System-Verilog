class axi_bfm;
	task run();
		$display("axi_bfm:: run");
	endtask
endclass
