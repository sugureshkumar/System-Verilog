library verilog;
use verilog.vl_types.all;
entity axi_tb is
end axi_tb;
