class axi_cov;
	task run();
		$display("axi_cov:: run");
	endtask
endclass
