program axi_tb;

	axi_env  env=new();
	initial begin
		env.run();
	end

endprogram
